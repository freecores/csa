// this key_schedule module
module key_schedule(i_ck,o_kk);
        input  [8*8-1:0]  i_ck;
        output [56*8-1:0] o_kk;

        wire   [64*8-1:0] kb;

        assign kb[(8*8)*8-1:(7*8)*8] = i_ck;

        key_perm k1( .i_key(kb[(8*8)*8-1:(7*8)*8]) ,.o_key(kb[(7*8)*8-1:(6*8)*8]));
        key_perm k2( .i_key(kb[(7*8)*8-1:(6*8)*8]) ,.o_key(kb[(6*8)*8-1:(5*8)*8]));
        key_perm k3( .i_key(kb[(6*8)*8-1:(5*8)*8]) ,.o_key(kb[(5*8)*8-1:(4*8)*8]));
        key_perm k4( .i_key(kb[(5*8)*8-1:(4*8)*8]) ,.o_key(kb[(4*8)*8-1:(3*8)*8]));
        key_perm k5( .i_key(kb[(4*8)*8-1:(3*8)*8]) ,.o_key(kb[(3*8)*8-1:(2*8)*8]));
        key_perm k6( .i_key(kb[(3*8)*8-1:(2*8)*8]) ,.o_key(kb[(2*8)*8-1:(1*8)*8]));
        key_perm k7( .i_key(kb[(2*8)*8-1:(1*8)*8]) ,.o_key(kb[(1*8)*8-1:(0*8)*8]));

        assign o_kk [(1*8)*8-1:(0*8)*8] = kb[(1*8)*8-1:(0*8)*8] ^ 64'h0000000000000000;
        assign o_kk [(2*8)*8-1:(1*8)*8] = kb[(2*8)*8-1:(1*8)*8] ^ 64'h0101010101010101;
        assign o_kk [(3*8)*8-1:(2*8)*8] = kb[(3*8)*8-1:(2*8)*8] ^ 64'h0202020202020202;
        assign o_kk [(4*8)*8-1:(3*8)*8] = kb[(4*8)*8-1:(3*8)*8] ^ 64'h0303030303030303;
        assign o_kk [(5*8)*8-1:(4*8)*8] = kb[(5*8)*8-1:(4*8)*8] ^ 64'h0404040404040404;
        assign o_kk [(6*8)*8-1:(5*8)*8] = kb[(6*8)*8-1:(5*8)*8] ^ 64'h0505050505050505;
        assign o_kk [(7*8)*8-1:(6*8)*8] = kb[(7*8)*8-1:(6*8)*8] ^ 64'h0606060606060606;

endmodule
