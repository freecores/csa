
// this module will do csa decrypt work
module decrypt(even_cw,odd_cw,encrypted,decrypted);
input  even_cw;
input  odd_cw;
input  encrypted;
output decrypted;

endmodule
